netcdf ww3.Point0_196806_spec {
dimensions:
	time = UNLIMITED ; // (55 currently)
	station = 1 ;
	string16 = 16 ;
	frequency = 24 ;
	direction = 24 ;
variables:
	double time(time) ;
		time:long_name = "julian day (UT)" ;
		time:standard_name = "time" ;
		time:calendar = "standard" ;
		time:units = "days since 1990-01-01 00:00:00" ;
		time:conventions = "Relative julian days with decimal part (as parts of the day)" ;
		time:axis = "T" ;
	int station(station) ;
		station:long_name = "station id" ;
		station:_FillValue = -2147483647 ;
		station:axis = "X" ;
	int string16(string16) ;
		string16:long_name = "station_name number of characters" ;
		string16:_FillValue = -2147483647 ;
		string16:axis = "W" ;
	char station_name(station, string16) ;
		station_name:long_name = "station name" ;
		station_name:content = "XW" ;
		station_name:associates = "station string16" ;
	float x(time, station) ;
		x:long_name = "x" ;
		x:standard_name = "x" ;
		x:globwave_name = "x" ;
		x:units = "m" ;
		x:scale_factor = 1.f ;
		x:add_offset = 0.f ;
		x:valid_min = 0.f ;
		x:valid_max = 10000.f ;
		x:_FillValue = 9.96921e+36f ;
		x:content = "TX" ;
		x:associates = "time station" ;
	float y(time, station) ;
		y:long_name = "y" ;
		y:standard_name = "y" ;
		y:globwave_name = "y" ;
		y:units = "m" ;
		y:scale_factor = 1.f ;
		y:add_offset = 0.f ;
		y:valid_min = 0.f ;
		y:valid_max = 10000.f ;
		y:_FillValue = 9.96921e+36f ;
		y:content = "TX" ;
		y:associates = "time station" ;
	float frequency(frequency) ;
		frequency:long_name = "frequency of center band" ;
		frequency:standard_name = "sea_surface_wave_frequency" ;
		frequency:globwave_name = "frequency" ;
		frequency:units = "s-1" ;
		frequency:scale_factor = 1.f ;
		frequency:add_offset = 0.f ;
		frequency:valid_min = 0.f ;
		frequency:valid_max = 10.f ;
		frequency:_FillValue = 9.96921e+36f ;
		frequency:axis = "Y" ;
	float frequency1(frequency) ;
		frequency1:long_name = "frequency of lower band" ;
		frequency1:standard_name = "frequency_of_lower_band" ;
		frequency1:globwave_name = "frequency_lower_band" ;
		frequency1:units = "s-1" ;
		frequency1:scale_factor = 1.f ;
		frequency1:add_offset = 0.f ;
		frequency1:valid_min = 0.f ;
		frequency1:valid_max = 10.f ;
		frequency1:_FillValue = 9.96921e+36f ;
		frequency1:content = "Y" ;
		frequency1:associates = "frequency" ;
	float frequency2(frequency) ;
		frequency2:long_name = "frequency of upper band" ;
		frequency2:standard_name = "frequency_of_upper_band" ;
		frequency2:globwave_name = "frequency_upper_band" ;
		frequency2:units = "s-1" ;
		frequency2:scale_factor = 1.f ;
		frequency2:add_offset = 0.f ;
		frequency2:valid_min = 0.f ;
		frequency2:valid_max = 10.f ;
		frequency2:_FillValue = 9.96921e+36f ;
		frequency2:content = "Y" ;
		frequency2:associates = "frequency" ;
	float direction(direction) ;
		direction:long_name = "sea surface wave to direction" ;
		direction:standard_name = "sea_surface_wave_to_direction" ;
		direction:globwave_name = "direction" ;
		direction:units = "degree" ;
		direction:scale_factor = 1.f ;
		direction:add_offset = 0.f ;
		direction:valid_min = 0.f ;
		direction:valid_max = 360.f ;
		direction:_FillValue = 9.96921e+36f ;
		direction:axis = "Z" ;
	float efth(time, station, frequency, direction) ;
		efth:long_name = "sea surface wave directional variance spectral density" ;
		efth:standard_name = "sea_surface_wave_directional_variance_spectral_density" ;
		efth:globwave_name = "directional_variance_spectral_density" ;
		efth:units = "m2 s rad-1" ;
		efth:scale_factor = 1.f ;
		efth:add_offset = 0.f ;
		efth:valid_min = 0.f ;
		efth:valid_max = 1.e+20f ;
		efth:_FillValue = 9.96921e+36f ;
		efth:content = "TXYZ" ;
		efth:associates = "time station frequency direction" ;
	float dpt(time, station) ;
		dpt:long_name = "depth" ;
		dpt:standard_name = "depth" ;
		dpt:globwave_name = "depth" ;
		dpt:units = "m" ;
		dpt:scale_factor = 1.f ;
		dpt:add_offset = 0.f ;
		dpt:valid_min = -100.f ;
		dpt:valid_max = 10000.f ;
		dpt:_FillValue = 9.96921e+36f ;
		dpt:content = "TX" ;
		dpt:associates = "time station" ;
	float wnd(time, station) ;
		wnd:long_name = "wind speed at 10m" ;
		wnd:standard_name = "wind_speed" ;
		wnd:globwave_name = "wind_speed" ;
		wnd:units = "m s-1" ;
		wnd:scale_factor = 1.f ;
		wnd:add_offset = 0.f ;
		wnd:valid_min = 0.f ;
		wnd:valid_max = 100.f ;
		wnd:_FillValue = 9.96921e+36f ;
		wnd:content = "TX" ;
		wnd:associates = "time station" ;
	float wnddir(time, station) ;
		wnddir:long_name = "wind direction" ;
		wnddir:standard_name = "wind_from_direction" ;
		wnddir:globwave_name = "wind_from_direction" ;
		wnddir:units = "degree" ;
		wnddir:scale_factor = 1.f ;
		wnddir:add_offset = 0.f ;
		wnddir:valid_min = 0.f ;
		wnddir:valid_max = 360.f ;
		wnddir:_FillValue = 9.96921e+36f ;
		wnddir:content = "TX" ;
		wnddir:associates = "time station" ;
	float cur(time, station) ;
		cur:long_name = "sea water speed" ;
		cur:standard_name = "sea_water_speed" ;
		cur:globwave_name = "sea_water_speed" ;
		cur:units = "m s-1" ;
		cur:scale_factor = 1.f ;
		cur:add_offset = 0.f ;
		cur:valid_min = 0.f ;
		cur:valid_max = 100.f ;
		cur:_FillValue = 9.96921e+36f ;
		cur:content = "TX" ;
		cur:associates = "time station" ;
	float curdir(time, station) ;
		curdir:long_name = "direction from of sea water velocity" ;
		curdir:standard_name = "direction_of_sea_water_velocity" ;
		curdir:globwave_name = "direction_of_sea_water_velocity" ;
		curdir:units = "degree" ;
		curdir:scale_factor = 1.f ;
		curdir:add_offset = 0.f ;
		curdir:valid_min = 0.f ;
		curdir:valid_max = 360.f ;
		curdir:_FillValue = 9.96921e+36f ;
		curdir:content = "TX" ;
		curdir:associates = "time station" ;

// global attributes:
		:product_name = "ww3.Point1_196806_spec.nc" ;
		:area = "1-D PROP. USING W3CSPC" ;
		:data_type = "OCO spectra 2D" ;
		:format_version = "1.1" ;
		:southernmost_latitude = "n/a" ;
		:northernmost_latitude = "n/a" ;
		:latitude_resolution = "n/a" ;
		:westernmost_longitude = "n/a" ;
		:easternmost_longitude = "n/a" ;
		:longitude_resolution = "n/a" ;
		:minimum_altitude = "n/a" ;
		:maximum_altitude = "n/a" ;
		:altitude_resolution = "n/a" ;
		:start_date = "1968-06-01 00:00:00" ;
		:stop_date = "1968-06-01 18:00:00" ;
		:field_type = "n/a" ;
data:

 time = -7884, -7883.98611111111, -7883.97222222222, -7883.95833333333, 
    -7883.94444444444, -7883.93055555556, -7883.91666666667, 
    -7883.90277777778, -7883.88888888889, -7883.875, -7883.86111111111, 
    -7883.84722222222, -7883.83333333333, -7883.81944444444, 
    -7883.80555555556, -7883.79166666667, -7883.77777777778, 
    -7883.76388888889, -7883.75, -7883.73611111111, -7883.72222222222, 
    -7883.70833333333, -7883.69444444444, -7883.68055555556, 
    -7883.66666666667, -7883.65277777778, -7883.63888888889, -7883.625, 
    -7883.61111111111, -7883.59722222222, -7883.58333333333, 
    -7883.56944444444, -7883.55555555556, -7883.54166666667, 
    -7883.52777777778, -7883.51388888889, -7883.5, -7883.48611111111, 
    -7883.47222222222, -7883.45833333333, -7883.44444444444, 
    -7883.43055555556, -7883.41666666667, -7883.40277777778, 
    -7883.38888888889, -7883.375, -7883.36111111111, -7883.34722222222, 
    -7883.33333333333, -7883.31944444444, -7883.30555555556, 
    -7883.29166666667, -7883.27777777778, -7883.26388888889, -7883.25 ;

 station = 1 ;

 string16 = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 station_name =
  "Point1" ;

 x =
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001,
  98.00001 ;

 y =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 frequency = 0.04, 0.044, 0.0484, 0.05324, 0.058564, 0.06442041, 0.07086245, 
    0.0779487, 0.08574356, 0.09431793, 0.1037497, 0.1141247, 0.1255372, 
    0.1380909, 0.1519, 0.16709, 0.183799, 0.2021789, 0.2223968, 0.2446365, 
    0.2691001, 0.2960101, 0.3256111, 0.3581723 ;

 frequency1 = 0.04, 0.042, 0.0462, 0.05082, 0.055902, 0.06149221, 0.06764143, 
    0.07440557, 0.08184613, 0.09003074, 0.09903383, 0.1089372, 0.1198309, 
    0.131814, 0.1449954, 0.159495, 0.1754445, 0.1929889, 0.2122878, 
    0.2335166, 0.2568683, 0.2825551, 0.3108106, 0.3418917 ;

 frequency2 = 0.042, 0.0462, 0.05082, 0.055902, 0.0614922, 0.06764143, 
    0.07440557, 0.08184613, 0.09003074, 0.09903383, 0.1089372, 0.1198309, 
    0.131814, 0.1449954, 0.159495, 0.1754445, 0.1929889, 0.2122878, 
    0.2335166, 0.2568683, 0.2825551, 0.3108106, 0.3418917, 0.3581723 ;

 direction = 90, 75, 60, 45, 30, 15, 0, 345, 330, 315, 300, 285, 270, 255, 
    240, 225, 210, 195, 180, 165, 150, 135, 120, 105 ;

 efth =
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604497, 0.521013, 0.2604497, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.000896766, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.000896766, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327485, 
    0.5616872, 1.12362, 0.5616872, 0.06327485, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255859e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255859e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116914e-07, 3.654561e-06, 7.310716e-06, 3.654561e-06, 4.116914e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 7.072087e-13, 3.70699e-07, 0.0003795956, 0.0218894, 
    0.1943109, 0.3887066, 0.1943109, 0.0218894, 0.0003795956, 3.70699e-07, 
    7.072087e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.175612e-13, 4.285427e-07, 0.0004388275, 0.02530501, 
    0.2246311, 0.4493602, 0.2246311, 0.02530501, 0.0004388275, 4.285427e-07, 
    8.175612e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.479257e-13, 4.968762e-07, 0.0005088008, 0.02934003, 
    0.2604498, 0.521013, 0.2604498, 0.02934003, 0.0005088008, 4.968762e-07, 
    9.479257e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.099978e-12, 5.765777e-07, 0.0005904153, 0.03404632, 
    0.3022272, 0.6045863, 0.3022272, 0.03404632, 0.0005904153, 5.765777e-07, 
    1.099978e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.273828e-12, 6.677049e-07, 0.0006837294, 0.03942729, 
    0.3499937, 0.7001401, 0.3499937, 0.03942729, 0.0006837294, 6.677049e-07, 
    1.273828e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.466641e-12, 7.687722e-07, 0.0007872221, 0.0453952, 
    0.4029705, 0.806117, 0.4029705, 0.0453952, 0.0007872221, 7.687722e-07, 
    1.466641e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.670727e-12, 8.757486e-07, 0.0008967661, 0.05171206, 
    0.4590449, 0.9182901, 0.4590449, 0.05171206, 0.0008967661, 8.757486e-07, 
    1.670727e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.871264e-12, 9.808646e-07, 0.001004405, 0.05791905, 
    0.514144, 1.028512, 0.514144, 0.05791905, 0.001004405, 9.808646e-07, 
    1.871264e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.044301e-12, 1.071566e-06, 0.001097283, 0.06327486, 
    0.5616872, 1.12362, 0.5616872, 0.06327486, 0.001097283, 1.071566e-06, 
    2.044301e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.156488e-12, 1.130371e-06, 0.001157499, 0.06674725, 
    0.5925114, 1.185281, 0.5925114, 0.06674725, 0.001157499, 1.130371e-06, 
    2.156488e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.168806e-12, 1.136827e-06, 0.00116411, 0.06712849, 
    0.5958956, 1.192051, 0.5958956, 0.06712849, 0.00116411, 1.136827e-06, 
    2.168806e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.046691e-12, 1.072819e-06, 0.001098566, 0.06334882, 
    0.5623438, 1.124933, 0.5623438, 0.06334882, 0.001098566, 1.072819e-06, 
    2.046691e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.77673e-12, 9.313122e-07, 0.0009536633, 0.05499304, 
    0.48817, 0.9765529, 0.48817, 0.05499304, 0.0009536633, 9.313122e-07, 
    1.77673e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.384251e-12, 7.255858e-07, 0.0007429995, 0.0428451, 
    0.3803335, 0.7608328, 0.3803335, 0.0428451, 0.0007429995, 7.255858e-07, 
    1.384251e-12, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 9.387728e-13, 4.920785e-07, 0.0005038881, 0.02905673, 
    0.2579349, 0.5159823, 0.2579349, 0.02905673, 0.0005038881, 4.920785e-07, 
    9.387728e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.336513e-13, 2.797251e-07, 0.0002864383, 0.01651748, 
    0.1466247, 0.2933134, 0.1466247, 0.01651748, 0.0002864383, 2.797251e-07, 
    5.336513e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.427098e-13, 1.272217e-07, 0.000130275, 0.007512312, 
    0.06668635, 0.1334018, 0.06668635, 0.007512312, 0.000130275, 
    1.272217e-07, 2.427098e-13, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 8.340111e-14, 4.371654e-08, 4.476571e-05, 0.002581417, 
    0.02291509, 0.04584017, 0.02291509, 0.002581417, 4.476571e-05, 
    4.371654e-08, 8.340111e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.018162e-14, 1.057864e-08, 1.083252e-05, 0.000624658, 
    0.005545052, 0.01109252, 0.005545052, 0.000624658, 1.083252e-05, 
    1.057864e-08, 2.018162e-14, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.154778e-15, 1.653646e-09, 1.693333e-06, 
    9.764611e-05, 0.0008667989, 0.001733976, 0.0008667989, 9.764611e-05, 
    1.693333e-06, 1.653646e-09, 3.154778e-15, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.866296e-16, 1.502432e-10, 1.53849e-07, 8.87171e-06, 
    7.875364e-05, 0.0001575417, 7.875364e-05, 8.87171e-06, 1.53849e-07, 
    1.502432e-10, 2.866296e-16, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.330104e-17, 6.972034e-12, 7.139358e-09, 
    4.116915e-07, 3.65456e-06, 7.310716e-06, 3.65456e-06, 4.116915e-07, 
    7.139358e-09, 6.972034e-12, 1.330104e-17, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 dpt =
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000,
  1000 ;

 wnd =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 wnddir =
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270 ;

 cur =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 curdir =
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270,
  270 ;
}
