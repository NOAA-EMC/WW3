netcdf ww3.Point1_196806_spec {
dimensions:
	time = UNLIMITED ; // (55 currently)
	station = 1 ;
	string40 = 40 ;
	frequency = 24 ;
	direction = 24 ;
variables:
	double time(time) ;
		time:long_name = "julian day (UT)" ;
		time:standard_name = "time" ;
		time:units = "days since 1990-01-01 00:00:00" ;
		time:conventions = "Relative julian days with decimal part (as parts of the day)" ;
		time:axis = "T" ;
		time:calendar = "standard" ;
	int station(station) ;
		station:long_name = "station id" ;
		station:_FillValue = -2147483647 ;
		station:axis = "X" ;
	int string40(string40) ;
		string40:long_name = "station_name number of characters" ;
		string40:_FillValue = -2147483647 ;
		string40:axis = "W" ;
	char station_name(station, string40) ;
		station_name:long_name = "station name" ;
		station_name:content = "XW" ;
		station_name:associates = "station string40" ;
	float x(time, station) ;
		x:long_name = "x" ;
		x:standard_name = "x" ;
		x:globwave_name = "x" ;
		x:units = "m" ;
		x:scale_factor = 1.f ;
		x:add_offset = 0.f ;
		x:valid_min = 0.f ;
		x:valid_max = 10000.f ;
		x:_FillValue = 9.96921e+36f ;
		x:content = "TX" ;
		x:associates = "time station" ;
	float y(time, station) ;
		y:long_name = "y" ;
		y:standard_name = "y" ;
		y:globwave_name = "y" ;
		y:units = "m" ;
		y:scale_factor = 1.f ;
		y:add_offset = 0.f ;
		y:valid_min = 0.f ;
		y:valid_max = 10000.f ;
		y:_FillValue = 9.96921e+36f ;
		y:content = "TX" ;
		y:associates = "time station" ;
	float frequency(frequency) ;
		frequency:long_name = "frequency of center band" ;
		frequency:standard_name = "sea_surface_wave_frequency" ;
		frequency:globwave_name = "frequency" ;
		frequency:units = "s-1" ;
		frequency:scale_factor = 1.f ;
		frequency:add_offset = 0.f ;
		frequency:valid_min = 0.f ;
		frequency:valid_max = 10.f ;
		frequency:_FillValue = 9.96921e+36f ;
		frequency:axis = "Y" ;
	float frequency1(frequency) ;
		frequency1:long_name = "frequency of lower band" ;
		frequency1:standard_name = "frequency_of_lower_band" ;
		frequency1:globwave_name = "frequency_lower_band" ;
		frequency1:units = "s-1" ;
		frequency1:scale_factor = 1.f ;
		frequency1:add_offset = 0.f ;
		frequency1:valid_min = 0.f ;
		frequency1:valid_max = 10.f ;
		frequency1:_FillValue = 9.96921e+36f ;
		frequency1:content = "Y" ;
		frequency1:associates = "frequency" ;
	float frequency2(frequency) ;
		frequency2:long_name = "frequency of upper band" ;
		frequency2:standard_name = "frequency_of_upper_band" ;
		frequency2:globwave_name = "frequency_upper_band" ;
		frequency2:units = "s-1" ;
		frequency2:scale_factor = 1.f ;
		frequency2:add_offset = 0.f ;
		frequency2:valid_min = 0.f ;
		frequency2:valid_max = 10.f ;
		frequency2:_FillValue = 9.96921e+36f ;
		frequency2:content = "Y" ;
		frequency2:associates = "frequency" ;
	float direction(direction) ;
		direction:long_name = "sea surface wave to direction" ;
		direction:standard_name = "sea_surface_wave_to_direction" ;
		direction:globwave_name = "direction" ;
		direction:units = "degree" ;
		direction:scale_factor = 1.f ;
		direction:add_offset = 0.f ;
		direction:valid_min = 0.f ;
		direction:valid_max = 360.f ;
		direction:_FillValue = 9.96921e+36f ;
		direction:axis = "Z" ;
	short efth(time, station, frequency, direction) ;
		efth:long_name = "sea surface wave directional variance spectral density" ;
		efth:globwave_name = "directional_variance_spectral_density" ;
		efth:standard_name = "base_ten_logarithm_of_sea_surface_wave_directional_variance_spectral_density" ;
		efth:units = "log10(m2 s rad-1 +1E-12)" ;
		efth:scale_factor = 0.0004f ;
		efth:add_offset = 0.f ;
		efth:valid_min = 0.f ;
		efth:valid_max = 1.e+20f ;
		efth:_FillValue = -32767s ;
		efth:content = "TXYZ" ;
		efth:associates = "time station frequency direction" ;
	short dpt(time, station) ;
		dpt:long_name = "depth" ;
		dpt:standard_name = "depth" ;
		dpt:globwave_name = "depth" ;
		dpt:units = "m" ;
		dpt:scale_factor = 0.5f ;
		dpt:add_offset = 0.f ;
		dpt:valid_min = -200 ;
		dpt:valid_max = 200000 ;
		dpt:_FillValue = -32767s ;
		dpt:content = "TX" ;
		dpt:associates = "time station" ;
	short wnd(time, station) ;
		wnd:long_name = "wind speed at 10m" ;
		wnd:standard_name = "wind_speed" ;
		wnd:globwave_name = "wind_speed" ;
		wnd:units = "m s-1" ;
		wnd:scale_factor = 0.1f ;
		wnd:add_offset = 0.f ;
		wnd:valid_min = 0 ;
		wnd:valid_max = 1000 ;
		wnd:_FillValue = -32767s ;
		wnd:content = "TX" ;
		wnd:associates = "time station" ;
	short wnddir(time, station) ;
		wnddir:long_name = "wind direction" ;
		wnddir:standard_name = "wind_from_direction" ;
		wnddir:globwave_name = "wind_from_direction" ;
		wnddir:units = "degree" ;
		wnddir:scale_factor = 0.1f ;
		wnddir:add_offset = 0.f ;
		wnddir:valid_min = 0 ;
		wnddir:valid_max = 3600 ;
		wnddir:_FillValue = -32767s ;
		wnddir:content = "TX" ;
		wnddir:associates = "time station" ;
	short cur(time, station) ;
		cur:long_name = "sea water speed" ;
		cur:standard_name = "sea_water_speed" ;
		cur:globwave_name = "sea_water_speed" ;
		cur:units = "m s-1" ;
		cur:scale_factor = 0.1f ;
		cur:add_offset = 0.f ;
		cur:valid_min = 0 ;
		cur:valid_max = 1000 ;
		cur:_FillValue = -32767s ;
		cur:content = "TX" ;
		cur:associates = "time station" ;
	short curdir(time, station) ;
		curdir:long_name = "direction from of sea water velocity" ;
		curdir:standard_name = "direction_of_sea_water_velocity" ;
		curdir:globwave_name = "direction_of_sea_water_velocity" ;
		curdir:units = "degree" ;
		curdir:scale_factor = 0.1f ;
		curdir:add_offset = 0.f ;
		curdir:valid_min = 0 ;
		curdir:valid_max = 3600 ;
		curdir:_FillValue = -32767s ;
		curdir:content = "TX" ;
		curdir:associates = "time station" ;

// global attributes:
		:product_name = "ww3.Point1_196806_spec.nc" ;
		:area = "1-D PROP. USING W3CSPC" ;
		:data_type = "OCO spectra 2D" ;
		:format_version = "1.1" ;
		:southernmost_latitude = "n/a" ;
		:northernmost_latitude = "n/a" ;
		:latitude_resolution = "n/a" ;
		:westernmost_longitude = "n/a" ;
		:easternmost_longitude = "n/a" ;
		:longitude_resolution = "n/a" ;
		:minimum_altitude = "n/a" ;
		:maximum_altitude = "n/a" ;
		:altitude_resolution = "n/a" ;
		:start_date = "1968-06-01 00:00:00" ;
		:stop_date = "1968-06-01 18:00:00" ;
		:field_type = "n/a" ;
data:

 time = -7884, -7883.98611111111, -7883.97222222222, -7883.95833333333, 
    -7883.94444444444, -7883.93055555556, -7883.91666666667, 
    -7883.90277777778, -7883.88888888889, -7883.875, -7883.86111111111, 
    -7883.84722222222, -7883.83333333333, -7883.81944444444, 
    -7883.80555555556, -7883.79166666667, -7883.77777777778, 
    -7883.76388888889, -7883.75, -7883.73611111111, -7883.72222222222, 
    -7883.70833333333, -7883.69444444444, -7883.68055555556, 
    -7883.66666666667, -7883.65277777778, -7883.63888888889, -7883.625, 
    -7883.61111111111, -7883.59722222222, -7883.58333333333, 
    -7883.56944444444, -7883.55555555556, -7883.54166666667, 
    -7883.52777777778, -7883.51388888889, -7883.5, -7883.48611111111, 
    -7883.47222222222, -7883.45833333333, -7883.44444444444, 
    -7883.43055555556, -7883.41666666667, -7883.40277777778, 
    -7883.38888888889, -7883.375, -7883.36111111111, -7883.34722222222, 
    -7883.33333333333, -7883.31944444444, -7883.30555555556, 
    -7883.29166666667, -7883.27777777778, -7883.26388888889, -7883.25 ;

 station = 1 ;

 string40 = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 station_name =
  "Point1" ;

 x =
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100,
  100 ;

 y =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 frequency = 0.04, 0.044, 0.0484, 0.05324, 0.058564, 0.06442041, 0.07086245, 
    0.0779487, 0.08574356, 0.09431793, 0.1037497, 0.1141247, 0.1255372, 
    0.1380909, 0.1519, 0.16709, 0.183799, 0.2021789, 0.2223968, 0.2446365, 
    0.2691001, 0.2960101, 0.3256111, 0.3581723 ;

 frequency1 = 0.04, 0.042, 0.0462, 0.05082, 0.055902, 0.06149221, 0.06764143, 
    0.07440557, 0.08184613, 0.09003074, 0.09903383, 0.1089372, 0.1198309, 
    0.131814, 0.1449954, 0.159495, 0.1754445, 0.1929889, 0.2122878, 
    0.2335166, 0.2568683, 0.2825551, 0.3108106, 0.3418917 ;

 frequency2 = 0.042, 0.0462, 0.05082, 0.055902, 0.0614922, 0.06764143, 
    0.07440557, 0.08184613, 0.09003074, 0.09903383, 0.1089372, 0.1198309, 
    0.131814, 0.1449954, 0.159495, 0.1754445, 0.1929889, 0.2122878, 
    0.2335166, 0.2568683, 0.2825551, 0.3108106, 0.3418917, 0.3581723 ;

 direction = 90, 75, 60, 45, 30, 15, 0, 345, 330, 315, 300, 285, 270, 255, 
    240, 225, 210, 195, 180, 165, 150, 135, 120, 105 ;

 efth =
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29419, -16077, 
    -8552, -4149, -1779, -1026, -1779, -4149, -8552, -16077, -29419, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29351, -15920, 
    -8394, -3992, -1621, -869, -1621, -3992, -8394, -15920, -29351, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29276, -15759, 
    -8234, -3831, -1461, -708, -1461, -3831, -8234, -15759, -29276, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29194, -15598, 
    -8072, -3670, -1299, -546, -1299, -3670, -8072, -15598, -29194, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29108, -15439, 
    -7913, -3511, -1140, -387, -1140, -3511, -7913, -15439, -29108, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29020, -15286, 
    -7760, -3357, -987, -234, -987, -3357, -7760, -15286, -29020, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28933, -15144, 
    -7618, -3216, -845, -93, -845, -3216, -7618, -15144, -28933, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28855, -15021, 
    -7495, -3093, -722, 31, -722, -3093, -7495, -15021, -28855, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28791, -14925, 
    -7399, -2997, -626, 127, -626, -2997, -7399, -14925, -28791, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28752, -14867, 
    -7341, -2939, -568, 185, -568, -2939, -7341, -14867, -28752, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28748, -14861, 
    -7335, -2933, -562, 191, -562, -2933, -7335, -14861, -28748, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28790, -14924, 
    -7398, -2996, -625, 128, -625, -2996, -7398, -14924, -28790, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -28891, -15077, 
    -7552, -3149, -779, -26, -779, -3149, -7552, -15077, -28891, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29057, -15348, 
    -7823, -3420, -1050, -297, -1050, -3420, -7823, -15348, -29057, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29281, -15770, 
    -8244, -3842, -1471, -718, -1471, -3842, -8244, -15770, -29281, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29536, -16383, 
    -8857, -4455, -2084, -1332, -2084, -4455, -8857, -16383, -29536, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29764, -17239, 
    -9713, -5311, -2940, -2187, -2940, -5311, -9713, -17239, -29764, -30000, 
    -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29913, -18398, 
    -10873, -6470, -4100, -3347, -4100, -6470, -10873, -18398, -29913, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29978, -19939, 
    -12413, -8011, -5640, -4887, -5640, -8011, -12413, -19939, -29978, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -29997, -21953, 
    -14428, -10026, -7655, -6902, -7655, -10026, -14428, -21953, -29997, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -24551, 
    -17032, -12630, -10259, -9507, -10259, -12630, -17032, -24551, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -27746, 
    -20366, -15964, -13593, -12840, -13593, -15964, -20366, -27746, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000,
  -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, -30000, 
    -30000, -30000, -30000, -30000, -30000, -30000 ;

 dpt =
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000,
  2000 ;

 wnd =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 wnddir =
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700 ;

 cur =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 curdir =
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700,
  2700 ;
}
